entity FA is
    port()